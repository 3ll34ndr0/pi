library ieee;

use ieee.std_logic_1164.all;

entity
  BrentKungFastAdder
is
port
  ( 
 
    
    a[0] : in std_logic
  ; a[1] : in std_logic
  ; a[2] : in std_logic
  ; a[3] : in std_logic
  ; b[0] : in std_logic
  ; b[1] : in std_logic
  ; b[2] : in std_logic
  ; b[3] : in std_logic

  
  ; sum[0] : out std_logic
  ; sum[1] : out std_logic
  ; sum[2] : out std_logic
  ; sum[3] : out std_logic
  ; cout : out std_logic
  );
end BrentKungFastAdder;

architecture
  structural
of
  BrentKungFastAdder
is
 --agregado para que Electric encuentre las celdas estandards
component and2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component or2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component xor2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component id
port( A : in std_logic;  Y : out std_logic);
 end component;
--
  signal w1 : std_logic;
  signal w2 : std_logic;
  signal w3 : std_logic;
  signal w4 : std_logic;
  signal w5 : std_logic;
  signal w6 : std_logic;
  signal w7 : std_logic;
  signal w8 : std_logic;
  signal w9 : std_logic;
  signal w10 : std_logic;
  signal w11 : std_logic;
  signal w12 : std_logic;
  signal w13 : std_logic;
  signal w14 : std_logic;
  signal w15 : std_logic;
  signal w16 : std_logic;
  signal w17 : std_logic;
  signal w18 : std_logic;
  signal w19 : std_logic;
  signal w20 : std_logic;
  signal w21 : std_logic;
  signal w22 : std_logic;
  signal w23 : std_logic;
  signal w24 : std_logic;
  signal w25 : std_logic;
  signal w26 : std_logic;
  signal w27 : std_logic;
  signal w28 : std_logic;
begin
-- deleted   c_w2      :  id    port map (a[0], a);
-- deleted   c_w3      :  id    port map (b[0], b);
  c_w1      :  xor2  port map (a, b, w1);
-- deleted   c_w6      :  id    port map (a[1], a);
-- deleted   c_w7      :  id    port map (b[1], b);
  c_w5      :  xor2  port map (a, b, w5);
  c_w8      :  and2  port map (a, b, w8);
  c_w4      :  xor2  port map (w5, w8, w4);
-- deleted   c_w11     :  id    port map (a[2], a);
-- deleted   c_w12     :  id    port map (b[2], b);
  c_w10     :  xor2  port map (a, b, w10);
  c_w14     :  and2  port map (a, b, w14);
  c_w15     :  and2  port map (w5, w8, w15);
  c_w13     :  or2   port map (w14, w15, w13);
  c_w9      :  xor2  port map (w10, w13, w9);
-- deleted   c_w18     :  id    port map (a[3], a);
-- deleted   c_w19     :  id    port map (b[3], b);
  c_w17     :  xor2  port map (a, b, w17);
  c_w21     :  and2  port map (a, b, w21);
  c_w22     :  and2  port map (w10, w13, w22);
  c_w20     :  or2   port map (w21, w22, w20);
  c_w16     :  xor2  port map (w17, w20, w16);
  c_w25     :  and2  port map (a, b, w25);
  c_w26     :  and2  port map (w17, w21, w26);
  c_w24     :  or2   port map (w25, w26, w24);
  c_w28     :  and2  port map (w17, w10, w28);
  c_w27     :  and2  port map (w28, w13, w27);
  c_w23     :  or2   port map (w24, w27, cout);

  
  c_sum[0]  :  id    port map (w1, sum[0]);
  c_sum[1]  :  id    port map (w4, sum[1]);
  c_sum[2]  :  id    port map (w9, sum[2]);
  c_sum[3]  :  id    port map (w16, sum[3]);
-- deleted --  c_cout    :  id    port map (cout, cout);
end structural;
