library ieee;

use ieee.std_logic_1164.all;

entity
  BrentKungFastAdder16
is
port
  ( 
 
    
    a[0] : in std_logic
  ; a[1] : in std_logic
  ; a[2] : in std_logic
  ; a[3] : in std_logic
  ; a[4] : in std_logic
  ; a[5] : in std_logic
  ; a[6] : in std_logic
  ; a[7] : in std_logic
  ; a[8] : in std_logic
  ; a[9] : in std_logic
  ; a[10] : in std_logic
  ; a[11] : in std_logic
  ; a[12] : in std_logic
  ; a[13] : in std_logic
  ; a[14] : in std_logic
  ; a[15] : in std_logic
  ; b[0] : in std_logic
  ; b[1] : in std_logic
  ; b[2] : in std_logic
  ; b[3] : in std_logic
  ; b[4] : in std_logic
  ; b[5] : in std_logic
  ; b[6] : in std_logic
  ; b[7] : in std_logic
  ; b[8] : in std_logic
  ; b[9] : in std_logic
  ; b[10] : in std_logic
  ; b[11] : in std_logic
  ; b[12] : in std_logic
  ; b[13] : in std_logic
  ; b[14] : in std_logic
  ; b[15] : in std_logic

  
  ; sum[0] : out std_logic
  ; sum[1] : out std_logic
  ; sum[2] : out std_logic
  ; sum[3] : out std_logic
  ; sum[4] : out std_logic
  ; sum[5] : out std_logic
  ; sum[6] : out std_logic
  ; sum[7] : out std_logic
  ; sum[8] : out std_logic
  ; sum[9] : out std_logic
  ; sum[10] : out std_logic
  ; sum[11] : out std_logic
  ; sum[12] : out std_logic
  ; sum[13] : out std_logic
  ; sum[14] : out std_logic
  ; sum[15] : out std_logic
  ; cout : out std_logic
  );
end BrentKungFastAdder16;

architecture
  structural
of
  BrentKungFastAdder16
is
 --agregado para que Electric encuentre las celdas estandards
component and2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component or2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component xor2
port( A, B : in std_logic;  Y : out std_logic);
 end component;
component id
port( A : in std_logic;  Y : out std_logic);
 end component;
--
  signal w1 : std_logic;
  signal w2 : std_logic;
  signal w3 : std_logic;
  signal w4 : std_logic;
  signal w5 : std_logic;
  signal w6 : std_logic;
  signal w7 : std_logic;
  signal w8 : std_logic;
  signal w9 : std_logic;
  signal w10 : std_logic;
  signal w11 : std_logic;
  signal w12 : std_logic;
  signal w13 : std_logic;
  signal w14 : std_logic;
  signal w15 : std_logic;
  signal w16 : std_logic;
  signal w17 : std_logic;
  signal w18 : std_logic;
  signal w19 : std_logic;
  signal w20 : std_logic;
  signal w21 : std_logic;
  signal w22 : std_logic;
  signal w23 : std_logic;
  signal w24 : std_logic;
  signal w25 : std_logic;
  signal w26 : std_logic;
  signal w27 : std_logic;
  signal w28 : std_logic;
  signal w29 : std_logic;
  signal w30 : std_logic;
  signal w31 : std_logic;
  signal w32 : std_logic;
  signal w33 : std_logic;
  signal w34 : std_logic;
  signal w35 : std_logic;
  signal w36 : std_logic;
  signal w37 : std_logic;
  signal w38 : std_logic;
  signal w39 : std_logic;
  signal w40 : std_logic;
  signal w41 : std_logic;
  signal w42 : std_logic;
  signal w43 : std_logic;
  signal w44 : std_logic;
  signal w45 : std_logic;
  signal w46 : std_logic;
  signal w47 : std_logic;
  signal w48 : std_logic;
  signal w49 : std_logic;
  signal w50 : std_logic;
  signal w51 : std_logic;
  signal w52 : std_logic;
  signal w53 : std_logic;
  signal w54 : std_logic;
  signal w55 : std_logic;
  signal w56 : std_logic;
  signal w57 : std_logic;
  signal w58 : std_logic;
  signal w59 : std_logic;
  signal w60 : std_logic;
  signal w61 : std_logic;
  signal w62 : std_logic;
  signal w63 : std_logic;
  signal w64 : std_logic;
  signal w65 : std_logic;
  signal w66 : std_logic;
  signal w67 : std_logic;
  signal w68 : std_logic;
  signal w69 : std_logic;
  signal w70 : std_logic;
  signal w71 : std_logic;
  signal w72 : std_logic;
  signal w73 : std_logic;
  signal w74 : std_logic;
  signal w75 : std_logic;
  signal w76 : std_logic;
  signal w77 : std_logic;
  signal w78 : std_logic;
  signal w79 : std_logic;
  signal w80 : std_logic;
  signal w81 : std_logic;
  signal w82 : std_logic;
  signal w83 : std_logic;
  signal w84 : std_logic;
  signal w85 : std_logic;
  signal w86 : std_logic;
  signal w87 : std_logic;
  signal w88 : std_logic;
  signal w89 : std_logic;
  signal w90 : std_logic;
  signal w91 : std_logic;
  signal w92 : std_logic;
  signal w93 : std_logic;
  signal w94 : std_logic;
  signal w95 : std_logic;
  signal w96 : std_logic;
  signal w97 : std_logic;
  signal w98 : std_logic;
  signal w99 : std_logic;
  signal w100 : std_logic;
  signal w101 : std_logic;
  signal w102 : std_logic;
  signal w103 : std_logic;
  signal w104 : std_logic;
  signal w105 : std_logic;
  signal w106 : std_logic;
  signal w107 : std_logic;
  signal w108 : std_logic;
  signal w109 : std_logic;
  signal w110 : std_logic;
  signal w111 : std_logic;
  signal w112 : std_logic;
  signal w113 : std_logic;
  signal w114 : std_logic;
  signal w115 : std_logic;
  signal w116 : std_logic;
  signal w117 : std_logic;
  signal w118 : std_logic;
  signal w119 : std_logic;
  signal w120 : std_logic;
  signal w121 : std_logic;
  signal w122 : std_logic;
  signal w123 : std_logic;
  signal w124 : std_logic;
  signal w125 : std_logic;
  signal w126 : std_logic;
  signal w127 : std_logic;
  signal w128 : std_logic;
  signal w129 : std_logic;
  signal w130 : std_logic;
  signal w131 : std_logic;
  signal w132 : std_logic;
  signal w133 : std_logic;
  signal w134 : std_logic;
  signal w135 : std_logic;
  signal w136 : std_logic;
  signal w137 : std_logic;
  signal w138 : std_logic;
  signal w139 : std_logic;
  signal w140 : std_logic;
  signal w141 : std_logic;
  signal w142 : std_logic;
begin
-- deleted   c_w2      :  id    port map (a[0], a);
-- deleted   c_w3      :  id    port map (b[0], b);
  c_w1      :  xor2  port map (a, b, w1);
-- deleted   c_w6      :  id    port map (a[1], a);
-- deleted   c_w7      :  id    port map (b[1], b);
  c_w5      :  xor2  port map (a, b, w5);
  c_w8      :  and2  port map (a, b, w8);
  c_w4      :  xor2  port map (w5, w8, w4);
-- deleted   c_w11     :  id    port map (a[2], a);
-- deleted   c_w12     :  id    port map (b[2], b);
  c_w10     :  xor2  port map (a, b, w10);
  c_w14     :  and2  port map (a, b, w14);
  c_w15     :  and2  port map (w5, w8, w15);
  c_w13     :  or2   port map (w14, w15, w13);
  c_w9      :  xor2  port map (w10, w13, w9);
-- deleted   c_w18     :  id    port map (a[3], a);
-- deleted   c_w19     :  id    port map (b[3], b);
  c_w17     :  xor2  port map (a, b, w17);
  c_w21     :  and2  port map (a, b, w21);
  c_w22     :  and2  port map (w10, w13, w22);
  c_w20     :  or2   port map (w21, w22, w20);
  c_w16     :  xor2  port map (w17, w20, w16);
-- deleted   c_w25     :  id    port map (a[4], a);
-- deleted   c_w26     :  id    port map (b[4], b);
  c_w24     :  xor2  port map (a, b, w24);
  c_w29     :  and2  port map (a, b, w29);
  c_w30     :  and2  port map (w17, w21, w30);
  c_w28     :  or2   port map (w29, w30, w28);
  c_w32     :  and2  port map (w17, w10, w32);
  c_w31     :  and2  port map (w32, w13, w31);
  c_w27     :  or2   port map (w28, w31, w27);
  c_w23     :  xor2  port map (w24, w27, w23);
-- deleted   c_w35     :  id    port map (a[5], a);
-- deleted   c_w36     :  id    port map (b[5], b);
  c_w34     :  xor2  port map (a, b, w34);
  c_w38     :  and2  port map (a, b, w38);
  c_w39     :  and2  port map (w24, w27, w39);
  c_w37     :  or2   port map (w38, w39, w37);
  c_w33     :  xor2  port map (w34, w37, w33);
-- deleted   c_w42     :  id    port map (a[6], a);
-- deleted   c_w43     :  id    port map (b[6], b);
  c_w41     :  xor2  port map (a, b, w41);
  c_w46     :  and2  port map (a, b, w46);
  c_w47     :  and2  port map (w34, w38, w47);
  c_w45     :  or2   port map (w46, w47, w45);
  c_w49     :  and2  port map (w34, w24, w49);
  c_w48     :  and2  port map (w49, w27, w48);
  c_w44     :  or2   port map (w45, w48, w44);
  c_w40     :  xor2  port map (w41, w44, w40);
-- deleted   c_w52     :  id    port map (a[7], a);
-- deleted   c_w53     :  id    port map (b[7], b);
  c_w51     :  xor2  port map (a, b, w51);
  c_w55     :  and2  port map (a, b, w55);
  c_w56     :  and2  port map (w41, w44, w56);
  c_w54     :  or2   port map (w55, w56, w54);
  c_w50     :  xor2  port map (w51, w54, w50);
-- deleted   c_w59     :  id    port map (a[8], a);
-- deleted   c_w60     :  id    port map (b[8], b);
  c_w58     :  xor2  port map (a, b, w58);
  c_w64     :  and2  port map (a, b, w64);
  c_w65     :  and2  port map (w51, w55, w65);
  c_w63     :  or2   port map (w64, w65, w63);
  c_w67     :  and2  port map (w51, w41, w67);
  c_w66     :  and2  port map (w67, w45, w66);
  c_w62     :  or2   port map (w63, w66, w62);
  c_w69     :  and2  port map (w67, w49, w69);
  c_w68     :  and2  port map (w69, w27, w68);
  c_w61     :  or2   port map (w62, w68, w61);
  c_w57     :  xor2  port map (w58, w61, w57);
-- deleted   c_w72     :  id    port map (a[9], a);
-- deleted   c_w73     :  id    port map (b[9], b);
  c_w71     :  xor2  port map (a, b, w71);
  c_w75     :  and2  port map (a, b, w75);
  c_w76     :  and2  port map (w58, w61, w76);
  c_w74     :  or2   port map (w75, w76, w74);
  c_w70     :  xor2  port map (w71, w74, w70);
-- deleted   c_w79     :  id    port map (a[10], a);
-- deleted   c_w80     :  id    port map (b[10], b);
  c_w78     :  xor2  port map (a, b, w78);
  c_w83     :  and2  port map (a, b, w83);
  c_w84     :  and2  port map (w71, w75, w84);
  c_w82     :  or2   port map (w83, w84, w82);
  c_w86     :  and2  port map (w71, w58, w86);
  c_w85     :  and2  port map (w86, w61, w85);
  c_w81     :  or2   port map (w82, w85, w81);
  c_w77     :  xor2  port map (w78, w81, w77);
-- deleted   c_w89     :  id    port map (a[11], a);
-- deleted   c_w90     :  id    port map (b[11], b);
  c_w88     :  xor2  port map (a, b, w88);
  c_w92     :  and2  port map (a, b, w92);
  c_w93     :  and2  port map (w78, w81, w93);
  c_w91     :  or2   port map (w92, w93, w91);
  c_w87     :  xor2  port map (w88, w91, w87);
-- deleted   c_w96     :  id    port map (a[12], a);
-- deleted   c_w97     :  id    port map (b[12], b);
  c_w95     :  xor2  port map (a, b, w95);
  c_w101    :  and2  port map (a, b, w101);
  c_w102    :  and2  port map (w88, w92, w102);
  c_w100    :  or2   port map (w101, w102, w100);
  c_w104    :  and2  port map (w88, w78, w104);
  c_w103    :  and2  port map (w104, w82, w103);
  c_w99     :  or2   port map (w100, w103, w99);
  c_w106    :  and2  port map (w104, w86, w106);
  c_w105    :  and2  port map (w106, w61, w105);
  c_w98     :  or2   port map (w99, w105, w98);
  c_w94     :  xor2  port map (w95, w98, w94);
-- deleted   c_w109    :  id    port map (a[13], a);
-- deleted   c_w110    :  id    port map (b[13], b);
  c_w108    :  xor2  port map (a, b, w108);
  c_w112    :  and2  port map (a, b, w112);
  c_w113    :  and2  port map (w95, w98, w113);
  c_w111    :  or2   port map (w112, w113, w111);
  c_w107    :  xor2  port map (w108, w111, w107);
-- deleted   c_w116    :  id    port map (a[14], a);
-- deleted   c_w117    :  id    port map (b[14], b);
  c_w115    :  xor2  port map (a, b, w115);
  c_w120    :  and2  port map (a, b, w120);
  c_w121    :  and2  port map (w108, w112, w121);
  c_w119    :  or2   port map (w120, w121, w119);
  c_w123    :  and2  port map (w108, w95, w123);
  c_w122    :  and2  port map (w123, w98, w122);
  c_w118    :  or2   port map (w119, w122, w118);
  c_w114    :  xor2  port map (w115, w118, w114);
-- deleted   c_w126    :  id    port map (a[15], a);
-- deleted   c_w127    :  id    port map (b[15], b);
  c_w125    :  xor2  port map (a, b, w125);
  c_w129    :  and2  port map (a, b, w129);
  c_w130    :  and2  port map (w115, w118, w130);
  c_w128    :  or2   port map (w129, w130, w128);
  c_w124    :  xor2  port map (w125, w128, w124);
  c_w135    :  and2  port map (a, b, w135);
  c_w136    :  and2  port map (w125, w129, w136);
  c_w134    :  or2   port map (w135, w136, w134);
  c_w138    :  and2  port map (w125, w115, w138);
  c_w137    :  and2  port map (w138, w119, w137);
  c_w133    :  or2   port map (w134, w137, w133);
  c_w140    :  and2  port map (w138, w123, w140);
  c_w139    :  and2  port map (w140, w99, w139);
  c_w132    :  or2   port map (w133, w139, w132);
  c_w142    :  and2  port map (w140, w106, w142);
  c_w141    :  and2  port map (w142, w61, w141);
  c_w131    :  or2   port map (w132, w141, cout);

  
  c_sum[0]  :  id    port map (w1, sum[0]);
  c_sum[1]  :  id    port map (w4, sum[1]);
  c_sum[2]  :  id    port map (w9, sum[2]);
  c_sum[3]  :  id    port map (w16, sum[3]);
  c_sum[4]  :  id    port map (w23, sum[4]);
  c_sum[5]  :  id    port map (w33, sum[5]);
  c_sum[6]  :  id    port map (w40, sum[6]);
  c_sum[7]  :  id    port map (w50, sum[7]);
  c_sum[8]  :  id    port map (w57, sum[8]);
  c_sum[9]  :  id    port map (w70, sum[9]);
  c_sum[10] :  id    port map (w77, sum[10]);
  c_sum[11] :  id    port map (w87, sum[11]);
  c_sum[12] :  id    port map (w94, sum[12]);
  c_sum[13] :  id    port map (w107, sum[13]);
  c_sum[14] :  id    port map (w114, sum[14]);
  c_sum[15] :  id    port map (w124, sum[15]);
-- deleted --  c_cout    :  id    port map (cout, cout);
end structural;
